VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

LAYER SVT_N
  TYPE IMPLANT ;
END SVT_N

LAYER GT
  TYPE MASTERSLICE ;
END GT

LAYER V0
  TYPE CUT ;
END V0

LAYER M1
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.096 ;
  WIDTH 0.032 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.032 WRONGDIRECTION ;" ;
END M1

LAYER V1
  TYPE CUT ;
END V1
LAYER M2
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION VERTICAL ;
  PITCH 0.052 ;
  WIDTH 0.024 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.024 WRONGDIRECTION ;" ;
END M2

LAYER V2
  TYPE CUT ;
END V2

LAYER M3
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.056 ;
  WIDTH 0.024 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.024 WRONGDIRECTION ;" ;
END M3

LAYER V3
  TYPE CUT ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.04 WRONGDIRECTION ;" ;
END M4
LAYER V4
  TYPE CUT ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.04 WRONGDIRECTION ;" ;
END M5

LAYER V5
  TYPE CUT ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.04 WRONGDIRECTION ;" ;
END M6

LAYER TV2
  TYPE CUT ;
END TV2

LAYER TM2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.72 ;
  WIDTH 0.36 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.36 WRONGDIRECTION ;" ;
END TM2
VIA V0
  LAYER GT ;
    RECT -0.021 -0.012 0.021 0.012 ;
  LAYER V0 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER M1 ;
    RECT -0.012 -0.048 0.012 0.048 ;
END V0

VIA V0_RH
  LAYER GT ;
    RECT -0.079 -0.016 0.079 0.016 ;
  LAYER V0 ;
    RECT -0.07 -0.016 0.07 0.016 ;
  LAYER M1 ;
    RECT -0.07 -0.052 0.07 0.052 ;
END V0_RH

VIA V0_RV
  LAYER GT ;
    RECT -0.025 -0.07 0.025 0.07 ;
  LAYER V0 ;
    RECT -0.016 -0.07 0.016 0.07 ;
  LAYER M1 ;
    RECT -0.016 -0.106 0.016 0.106 ;
END V0_RV
SITE 96s6t_CoreSite
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.096 BY 0.384 ;
END 96s6t_CoreSite

MACRO OR2V1_96S6T24UL
  CLASS CORE ;
  FOREIGN OR2V1_96S6T24UL ;
  ORIGIN 0 0 ;
  SIZE 0.384 BY 0.384 ;
  SYMMETRY X Y ;
  SITE 96s6t_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.06 0.166 0.092 0.198 ;
      LAYER M1 ;
        RECT 0.029 0.112 0.101 0.222 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.17 0.176 0.202 0.208 ;
      LAYER M1 ;
        RECT 0.159 0.112 0.211 0.272 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V0 ;
        RECT -0.016 0.368 0.016 0.4 ;
        RECT 0.08 0.368 0.112 0.4 ;
        RECT 0.176 0.368 0.208 0.4 ;
        RECT 0.272 0.368 0.304 0.4 ;
        RECT 0.368 0.368 0.4 0.4 ;
      LAYER M1 ;
        RECT -0.048 0.368 0.432 0.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V0 ;
        RECT -0.016 -0.016 0.016 0.016 ;
        RECT 0.08 -0.016 0.112 0.016 ;
        RECT 0.176 -0.016 0.208 0.016 ;
        RECT 0.272 -0.016 0.304 0.016 ;
        RECT 0.368 -0.016 0.4 0.016 ;
      LAYER M1 ;
        RECT -0.048 -0.016 0.432 0.016 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.32 0.099 0.352 0.131 ;
        RECT 0.32 0.253 0.352 0.285 ;
      LAYER M1 ;
        POLYGON 0.353 0.31 0.353 0.074 0.307 0.074 0.307 0.12 0.316 0.12 0.316 0.264 0.307 0.264 0.307 0.31 ;
    END
    ANTENNADIFFAREA 0.016128 ;
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.096 -0.096 0.48 0.192 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.096 0.192 0.48 0.48 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      POLYGON 0.275 0.336 0.275 0.24 0.283 0.24 0.283 0.144 0.275 0.144 0.275 0.048 0.103 0.048 0.103 0.08 0.243 0.08 0.243 0.304 0.076 0.304 0.076 0.254 0.029 0.254 0.029 0.336 ;
    LAYER AA ;
      RECT 0 0.24 0.384 0.336 ;
      RECT 0 0.048 0.384 0.144 ;
    LAYER ULVT_N ;
      RECT 0 0 0.384 0.192 ;
    LAYER ULVT_P ;
      RECT 0 0.192 0.384 0.384 ;
  END
END OR2V1_96S6T24UL

MACRO AND2V1_96S6T24UL
  CLASS CORE ;
  FOREIGN AND2V1_96S6T24UL ;
  ORIGIN 0 0 ;
  SIZE 0.384 BY 0.384 ;
  SYMMETRY X Y ;
  SITE 96s6t_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.06 0.186 0.092 0.218 ;
      LAYER M1 ;
        RECT 0.029 0.162 0.101 0.272 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.17 0.176 0.202 0.208 ;
      LAYER M1 ;
        RECT 0.159 0.112 0.211 0.272 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V0 ;
        RECT -0.016 0.368 0.016 0.4 ;
        RECT 0.08 0.368 0.112 0.4 ;
        RECT 0.176 0.368 0.208 0.4 ;
        RECT 0.272 0.368 0.304 0.4 ;
        RECT 0.368 0.368 0.4 0.4 ;
      LAYER M1 ;
        RECT -0.048 0.368 0.432 0.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V0 ;
        RECT -0.016 -0.016 0.016 0.016 ;
        RECT 0.08 -0.016 0.112 0.016 ;
        RECT 0.176 -0.016 0.208 0.016 ;
        RECT 0.272 -0.016 0.304 0.016 ;
        RECT 0.368 -0.016 0.4 0.016 ;
      LAYER M1 ;
        RECT -0.048 -0.016 0.432 0.016 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.32 0.099 0.352 0.131 ;
        RECT 0.32 0.253 0.352 0.285 ;
      LAYER M1 ;
        POLYGON 0.353 0.31 0.353 0.074 0.307 0.074 0.307 0.12 0.316 0.12 0.316 0.264 0.307 0.264 0.307 0.31 ;
    END
    ANTENNADIFFAREA 0.016128 ;
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.096 -0.096 0.48 0.192 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      POLYGON 0.275 0.336 0.275 0.24 0.283 0.24 0.283 0.144 0.275 0.144 0.275 0.048 0.029 0.048 0.029 0.13 0.076 0.13 0.076 0.08 0.243 0.08 0.243 0.304 0.103 0.304 0.103 0.336 ;
    LAYER AA ;
      RECT 0 0.24 0.384 0.336 ;
      RECT 0 0.048 0.384 0.144 ;
    LAYER ULVT_N ;
      RECT 0 0 0.384 0.192 ;
    LAYER ULVT_P ;
      RECT 0 0.192 0.384 0.384 ;
  END
END AND2V1_96S6T24UL

MACRO CLKINV1_96S6T24UL
  CLASS CORE ;
  FOREIGN CLKINV1_96S6T24UL ;
  ORIGIN 0 0 ;
  SIZE 0.192 BY 0.384 ;
  SYMMETRY X Y ;
  SITE 96s6t_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.052 0.176 0.084 0.208 ;
      LAYER M1 ;
        RECT 0.038 0.1 0.091 0.284 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V0 ;
        RECT -0.016 0.368 0.016 0.4 ;
        RECT 0.08 0.368 0.112 0.4 ;
        RECT 0.176 0.368 0.208 0.4 ;
      LAYER M1 ;
        RECT -0.048 0.368 0.24 0.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V0 ;
        RECT -0.016 -0.016 0.016 0.016 ;
        RECT 0.08 -0.016 0.112 0.016 ;
        RECT 0.176 -0.016 0.208 0.016 ;
      LAYER M1 ;
        RECT -0.048 -0.016 0.24 0.016 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.128 0.088 0.16 0.12 ;
        RECT 0.128 0.264 0.16 0.296 ;
      LAYER M1 ;
        RECT 0.125 0.056 0.163 0.328 ;
    END
    ANTENNADIFFAREA 0.016128 ;
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.096 -0.096 0.288 0.192 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.096 0.192 0.288 0.48 ;
    END
  END VNW
  OBS
    LAYER AA ;
      RECT 0 0.24 0.192 0.336 ;
      RECT 0 0.048 0.192 0.144 ;
    LAYER ULVT_N ;
      RECT 0 0 0.192 0.192 ;
    LAYER ULVT_P ;
      RECT 0 0.192 0.192 0.384 ;
  END
END CLKINV1_96S6T24UL
MACRO CLKNAND2V1_96S6T24UL
  CLASS CORE ;
  FOREIGN CLKNAND2V1_96S6T24UL ;
  ORIGIN 0 0 ;
  SIZE 0.288 BY 0.384 ;
  SYMMETRY X Y ;
  SITE 96s6t_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.152 0.176 0.184 0.208 ;
      LAYER M1 ;
        RECT 0.136 0.1 0.19 0.266 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.052 0.176 0.084 0.208 ;
      LAYER M1 ;
        RECT 0.04 0.056 0.086 0.233 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V0 ;
        RECT -0.016 0.368 0.016 0.4 ;
        RECT 0.08 0.368 0.112 0.4 ;
        RECT 0.176 0.368 0.208 0.4 ;
        RECT 0.272 0.368 0.304 0.4 ;
      LAYER M1 ;
        RECT -0.048 0.368 0.336 0.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V0 ;
        RECT -0.016 -0.016 0.016 0.016 ;
        RECT 0.08 -0.016 0.112 0.016 ;
        RECT 0.176 -0.016 0.208 0.016 ;
        RECT 0.272 -0.016 0.304 0.016 ;
      LAYER M1 ;
        RECT -0.048 -0.016 0.336 0.016 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.224 0.097 0.256 0.129 ;
        RECT 0.128 0.304 0.16 0.336 ;
      LAYER M1 ;
        POLYGON 0.259 0.336 0.259 0.072 0.222 0.072 0.222 0.299 0.092 0.299 0.092 0.336 ;
    END
    ANTENNADIFFAREA 0.014976 ;
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.096 -0.096 0.384 0.192 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.096 0.192 0.384 0.48 ;
    END
  END VNW
  OBS
    LAYER AA ;
      RECT 0 0.24 0.288 0.336 ;
      RECT 0 0.048 0.288 0.144 ;
    LAYER ULVT_N ;
      RECT 0 0 0.288 0.192 ;
    LAYER ULVT_P ;
      RECT 0 0.192 0.288 0.384 ;
  END
END CLKNAND2V1_96S6T24UL

MACRO NAND2BV1_96S6T24UL
  CLASS CORE ;
  FOREIGN NAND2BV1_96S6T24UL ;
  ORIGIN 0 0 ;
  SIZE 0.384 BY 0.384 ;
  SYMMETRY X Y ;
  SITE 96s6t_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER V0 ;
        RECT -0.016 0.368 0.016 0.4 ;
        RECT 0.08 0.368 0.112 0.4 ;
        RECT 0.176 0.368 0.208 0.4 ;
        RECT 0.272 0.368 0.304 0.4 ;
        RECT 0.368 0.368 0.4 0.4 ;
      LAYER M1 ;
        RECT -0.048 0.368 0.432 0.4 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER V0 ;
        RECT -0.016 -0.016 0.016 0.016 ;
        RECT 0.08 -0.016 0.112 0.016 ;
        RECT 0.176 -0.016 0.208 0.016 ;
        RECT 0.272 -0.016 0.304 0.016 ;
        RECT 0.368 -0.016 0.4 0.016 ;
      LAYER M1 ;
        RECT -0.048 -0.016 0.432 0.016 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.032 0.081 0.064 0.113 ;
        RECT 0.128 0.304 0.16 0.336 ;
      LAYER M1 ;
        POLYGON 0.185 0.336 0.185 0.304 0.066 0.304 0.066 0.056 0.029 0.056 0.029 0.336 ;
    END
    ANTENNADIFFAREA 0.014976 ;
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.254 0.183 0.286 0.215 ;
      LAYER V1 ;
        RECT 0.262 0.232 0.286 0.256 ;
      LAYER M2 ;
        RECT 0.122 0.232 0.322 0.256 ;
    END
    ANTENNAPARTIALMETALAREA 0.005143 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER TM2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER ALPA ;
    ANTENNAPARTIALCUTAREA 0.000576 LAYER V1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
    ANTENNAMAXAREACAR 1.116102 LAYER M1 ;
    ANTENNAMAXAREACAR 1.116102 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER TM2 ;
    ANTENNAMAXAREACAR 0 LAYER ALPA ;
    ANTENNAMAXCUTCAR 0.125 LAYER V1 ;
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER V0 ;
        RECT 0.177 0.161 0.209 0.193 ;
      LAYER V1 ;
        RECT 0.167 0.18 0.191 0.204 ;
      LAYER M2 ;
        RECT 0.107 0.18 0.307 0.204 ;
    END
    ANTENNAPARTIALMETALAREA 0.005184 LAYER M1 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER TM2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER ALPA ;
    ANTENNAPARTIALCUTAREA 0.000576 LAYER V1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.004608 ;
    ANTENNAMAXAREACAR 1.125 LAYER M1 ;
    ANTENNAMAXAREACAR 1.125 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER TM2 ;
    ANTENNAMAXAREACAR 0 LAYER ALPA ;
    ANTENNAMAXCUTCAR 0.125 LAYER V1 ;
  END B1
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.096 -0.096 0.48 0.192 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.096 0.192 0.48 0.48 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      POLYGON 0.355 0.31 0.355 0.054 0.266 0.054 0.266 0.1 0.318 0.1 0.318 0.31 ;
      RECT 0.249 0.14 0.286 0.279 ;
      RECT 0.167 0.138 0.215 0.246 ;
      POLYGON 0.135 0.242 0.135 0.106 0.182 0.106 0.182 0.074 0.098 0.074 0.098 0.242 ;
    LAYER M2 ;
      RECT 0.101 0.076 0.348 0.1 ;
    LAYER V1 ;
      RECT 0.291 0.076 0.315 0.1 ;
      RECT 0.133 0.076 0.157 0.1 ;
    LAYER AA ;
      RECT 0 0.24 0.384 0.336 ;
      RECT 0 0.048 0.384 0.144 ;
    LAYER ULVT_N ;
      RECT 0 0 0.384 0.192 ;
    LAYER ULVT_P ;
      RECT 0 0.192 0.384 0.384 ;
  END
END NAND2BV1_96S6T24UL

END LIBRARY

